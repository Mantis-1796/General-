module dut(input clk,rst,)
