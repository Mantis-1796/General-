TYPE : 1
module half_adder(input wire clk,
                  input wire rst,
                  input wire a,
                  input wire b,
                  output reg sum);
TYPE : 2
module half_adder(input clk,
                  input rst,
                  input a,
                  input b,
                  output reg sum);
TYPE : 3
module half_adder(clk,rst,a,b,sum);
    input clk;
    input rst;
    input a,b;
    output reg sum;
